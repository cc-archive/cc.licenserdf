<!DOCTYPE html PUBLIC "-//W3C//DTD XHTML+RDFa 1.0//EN" "http://www.w3.org/MarkUp/DTD/xhtml-rdfa-1.dtd">
<html xmlns="http://www.w3.org/1999/xhtml"
      xmlns:cc="http://creativecommons.org/ns#"
      xmlns:dc="http://purl.org/dc/elements/1.1/">
  <head>
    <title>Creative Commons &mdash;
      Erkännande 3.0 Hong Kong
    </title><link rel="stylesheet" type="text/css" href="http://yui.yahooapis.com/2.6.0/build/container/assets/skins/sam/container.css" /> 

    <link rel="stylesheet" type="text/css"
          href="http://creativecommons.org/@@/cc/includes/deed3.css"
          media="screen" />
    
    <link rel="stylesheet" type="text/css"
          href="http://creativecommons.org/@@/cc/includes/deed3-print.css"
          media="print" />
    <link rel="stylesheet" type="text/css"
          href="http://creativecommons.org/@@/cc/includes/jurisdictions.css"
          media="screen" />

    <!--[if lt IE 7]><link rel="stylesheet" type="text/css" href="/includes/deed3-ie.css" media="screen" tal:attributes="href context/++resource++cc/includes/deed3-ie.css" /><![endif]-->

    <link rel="alternate" type="application/rdf+xml" href="rdf" /> 
    

<script type="text/javascript">
function setCookie(name, value, expires, path, domain, secure) {
    document.cookie= name + "=" + escape(value) +
        ((expires) ? "; expires=" + expires.toGMTString() : "") +
        ((path) ? "; path=" + path : "") +
        ((domain) ? "; domain=" + domain : "") +
        ((secure) ? "; secure" : "");
}
var expiry = new Date();
expiry.setTime(expiry.getTime()+(5*365*24*60*60*1000));
setCookie('lang','%s', expiry, '/');
</script>



    <script type="text/javascript" src="http://yui.yahooapis.com/2.6.0/build/yahoo-dom-event/yahoo-dom-event.js">
    </script> 
    <script type="text/javascript" src="http://yui.yahooapis.com/2.6.0/build/connection/connection-min.js">
    </script> 
    <script type="text/javascript" src="http://yui.yahooapis.com/2.6.0/build/json/json-min.js">
    </script>

    <script type="text/javascript"
            src="http://creativecommons.org/@@/cc/includes/referrer/deed.js">
    </script>

    <script type="text/javascript" src="http://yui.yahooapis.com/2.6.0/build/container/container-min.js">
    </script>

    <script type="text/javascript"
            src="http://creativecommons.org/@@/cc/includes/help.js">
    </script>

    <script src="http://www.google-analytics.com/urchin.js" type="text/javascript"></script>
    <script type="text/javascript">
        _uacct="UA-2010376-1";  urchinTracker();
    </script>

   

  </head>
  <body class="yui-skin-sam">

    <!-- 
<rdf:RDF xmlns="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <License rdf:about="http://creativecommons.org/licenses/by/3.0/hk/">
        <permits rdf:resource="http://creativecommons.org/ns#Reproduction"/>
        <permits rdf:resource="http://creativecommons.org/ns#Distribution"/>
        <requires rdf:resource="http://creativecommons.org/ns#Notice"/>
        <requires rdf:resource="http://creativecommons.org/ns#Attribution"/>
        <permits rdf:resource="http://creativecommons.org/ns#DerivativeWorks"/>
      </License>
    </rdf:RDF>
   -->

    <div id="header">

    

<div id="languages">
<span style="text-align:left" dir="ltr">Denna sida finns tillgänglig på följande språk:</span>
<br />



<a href="./deed.af" title="Afrikaans" hreflang="af"
   rel="alternate nofollow" xml:lang="af">Afrikaans</a>




<a href="./deed.bg" title="български" hreflang="bg"
   rel="alternate nofollow" xml:lang="bg">български</a>




<a href="./deed.ca" title="Català" hreflang="ca"
   rel="alternate nofollow" xml:lang="ca">Català</a>




<a href="./deed.cs" title="Česko" hreflang="cs"
   rel="alternate nofollow" xml:lang="cs">Česko</a>




<a href="./deed.da" title="Dansk" hreflang="da"
   rel="alternate nofollow" xml:lang="da">Dansk</a>




<a href="./deed.de" title="Deutsch" hreflang="de"
   rel="alternate nofollow" xml:lang="de">Deutsch</a>




<a href="./deed.en" title="English" hreflang="en"
   rel="alternate nofollow" xml:lang="en">English</a>




<a href="./deed.en_CA" title="English (CA)" hreflang="en_CA"
   rel="alternate nofollow" xml:lang="en_CA">English (CA)</a>




<a href="./deed.en_GB" title="English (GB)" hreflang="en_GB"
   rel="alternate nofollow" xml:lang="en_GB">English (GB)</a>




<a href="./deed.en_HK" title="English (Hong Kong)"
   hreflang="en_HK" rel="alternate nofollow"
   xml:lang="en_HK">English (Hong Kong)</a>




<a href="./deed.en_SG" title="English (Singapore)"
   hreflang="en_SG" rel="alternate nofollow"
   xml:lang="en_SG">English (Singapore)</a>




<a href="./deed.en_US" title="English (US)" hreflang="en_US"
   rel="alternate nofollow" xml:lang="en_US">English (US)</a>




<a href="./deed.eo" title="Esperanto" hreflang="eo"
   rel="alternate nofollow" xml:lang="eo">Esperanto</a>




<a href="./deed.es" title="Castellano" hreflang="es"
   rel="alternate nofollow" xml:lang="es">Castellano</a>




<a href="./deed.es_AR" title="Castellano (AR)"
   hreflang="es_AR" rel="alternate nofollow"
   xml:lang="es_AR">Castellano (AR)</a>




<a href="./deed.es_CL" title="Español (CL)" hreflang="es_CL"
   rel="alternate nofollow" xml:lang="es_CL">Español (CL)</a>




<a href="./deed.es_CO" title="Castellano (CO)"
   hreflang="es_CO" rel="alternate nofollow"
   xml:lang="es_CO">Castellano (CO)</a>




<a href="./deed.es_EC" title="Español (Ecuador)"
   hreflang="es_EC" rel="alternate nofollow"
   xml:lang="es_EC">Español (Ecuador)</a>




<a href="./deed.es_GT" title="Español (Guatemala)"
   hreflang="es_GT" rel="alternate nofollow"
   xml:lang="es_GT">Español (Guatemala)</a>




<a href="./deed.es_MX" title="Castellano (MX)"
   hreflang="es_MX" rel="alternate nofollow"
   xml:lang="es_MX">Castellano (MX)</a>




<a href="./deed.es_PE" title="Castellano (PE)"
   hreflang="es_PE" rel="alternate nofollow"
   xml:lang="es_PE">Castellano (PE)</a>




<a href="./deed.eu" title="Euskara" hreflang="eu"
   rel="alternate nofollow" xml:lang="eu">Euskara</a>




<a href="./deed.fi" title="Suomeksi" hreflang="fi"
   rel="alternate nofollow" xml:lang="fi">Suomeksi</a>




<a href="./deed.fr" title="français" hreflang="fr"
   rel="alternate nofollow" xml:lang="fr">français</a>




<a href="./deed.fr_CA" title="français (CA)"
   hreflang="fr_CA" rel="alternate nofollow"
   xml:lang="fr_CA">français (CA)</a>




<a href="./deed.gl" title="Galego" hreflang="gl"
   rel="alternate nofollow" xml:lang="gl">Galego</a>




<a href="./deed.he" title="עברית" hreflang="he"
   rel="alternate nofollow" xml:lang="he">עברית</a>




<a href="./deed.hr" title="hrvatski" hreflang="hr"
   rel="alternate nofollow" xml:lang="hr">hrvatski</a>




<a href="./deed.hu" title="Magyar" hreflang="hu"
   rel="alternate nofollow" xml:lang="hu">Magyar</a>




<a href="./deed.it" title="Italiano" hreflang="it"
   rel="alternate nofollow" xml:lang="it">Italiano</a>




<a href="./deed.ja" title="日本語" hreflang="ja"
   rel="alternate nofollow" xml:lang="ja">日本語</a>




<a href="./deed.ko" title="한국어" hreflang="ko"
   rel="alternate nofollow" xml:lang="ko">한국어</a>




<a href="./deed.mk" title="Macedonian" hreflang="mk"
   rel="alternate nofollow" xml:lang="mk">Macedonian</a>




<a href="./deed.ms" title="Melayu" hreflang="ms"
   rel="alternate nofollow" xml:lang="ms">Melayu</a>




<a href="./deed.nl" title="Nederlands" hreflang="nl"
   rel="alternate nofollow" xml:lang="nl">Nederlands</a>




<a href="./deed.no" title="Norsk" hreflang="no"
   rel="alternate nofollow" xml:lang="no">Norsk</a>




<a href="./deed.nso" title="Sesotho sa Leboa" hreflang="nso"
   rel="alternate nofollow" xml:lang="nso">Sesotho sa Leboa</a>




<a href="./deed.pl" title="polski" hreflang="pl"
   rel="alternate nofollow" xml:lang="pl">polski</a>




<a href="./deed.pt" title="Português" hreflang="pt"
   rel="alternate nofollow" xml:lang="pt">Português</a>




<a href="./deed.ro" title="română" hreflang="ro"
   rel="alternate nofollow" xml:lang="ro">română</a>




<a href="./deed.sl" title="slovenski jezik" hreflang="sl"
   rel="alternate nofollow" xml:lang="sl">slovenski jezik</a>




<a href="./deed.sr" title="српски " hreflang="sr"
   rel="alternate nofollow" xml:lang="sr">српски </a>




<a href="./deed.sr_LATN" title="srpski (latinica)"
   hreflang="sr_LATN" rel="alternate nofollow"
   xml:lang="sr_LATN">srpski (latinica)</a>




<a href="./deed.st" title="Sotho" hreflang="st"
   rel="alternate nofollow" xml:lang="st">Sotho</a>




<a href="./deed.sv" title="svenska" hreflang="sv"
   rel="alternate nofollow" xml:lang="sv">svenska</a>




<a href="./deed.th" title="ไทย" hreflang="th"
   rel="alternate nofollow" xml:lang="th">ไทย</a>




<a href="./deed.zh" title="中文" hreflang="zh"
   rel="alternate nofollow" xml:lang="zh">中文</a>




<a href="./deed.zh_HK" title="中文（香港）" hreflang="zh_HK"
   rel="alternate nofollow" xml:lang="zh_HK">中文（香港）</a>




<a href="./deed.zh_TW" title="華語 (台灣)" hreflang="zh_TW"
   rel="alternate nofollow" xml:lang="zh_TW">華語 (台灣)</a>




<a href="./deed.zu" title="isiZulu" hreflang="zu"
   rel="alternate nofollow" xml:lang="zu">isiZulu</a>


</div>


    </div>

    <div id="deed" style="text-align:left" class="green"
         dir="ltr">

      <div id="deed-head">
	<div id="cc-logo">
	  <img src="/images/deed/cc-logo.jpg" alt="cc logo">
	</div>
	<div id="cc-link">
	  <a rel="dc:creator" href="http://creativecommons.org/">
            <span property="dc:title">Creative Commons</span>
          </a>	       
	</div>
	<h1><span>Creative Commons License Deed</span></h1>

        <div id="deed-license">
	        <h2 property="dc:title">Erkännande 3.0 Hong Kong</h2>
        </div>
      </div>

      <div id="deed-main" style="text-align:left" dir="ltr">
       <div id="deed-main-content" class="hk">

          
  <div id="libre">
    <a href="http://freedomdefined.org/">
      <img src="/images/deed/seal.png" style="border: 0"
           alt="This license is acceptable for Free Cultural Works." />
    </a>
  </div>

        <div id="deed-rights" style="text-align:left"
             dir="ltr">

        

<a href="/worldwide/hk/"><img
    src="/images/international/hk.png" style="border: 0"
    alt="hk" /></a>
<h3 rel="cc:permits"
    resource="http://creativecommons.org/ns#Reproduction">Du får:</h3>
		      <ul class="license-properties">
			<li class="license share" rel="cc:permits"
       resource="http://creativecommons.org/ns#Distribution"><strong>att Dela</strong> — att kopiera, distribuera och sända verket</li>
			      <li class="license remix" rel="cc:permits"
             resource="http://creativecommons.org/ns#DerivativeWorks"><strong>att Remixa</strong> — att skapa bearbetningar</li>
            <li id="more-container" class="license-hidden"><span id="devnations-container" /></li>
		      </ul>
        </div>
        <div id="deed-conditions">
	  <h3>På följande villkor:</h3>

	  <ul class="license-properties" style="text-align:left"
       dir="ltr"> 
            <li rel="cc:requires"
                resource="http://creativecommons.org/ns#Attribution"
                class="license by">
	      <p><strong>Erkännande</strong> &mdash;
		<span id="attribution-container">Du måste ange upphovsmannen och/eller licensgivaren på det sätt de anger (men inte på ett sätt som antyder att de godkänt eller rekommenderar din använding av verket).</span>
		
		<span id="by-more-container" />
	      </p>

	      
		<p id="work-attribution-container" style="display:none;">
		  <strong>Attribute this work:</strong><br />
		  <input id="work-attribution" value="" type="text" readonly="readonly" onclick="this.select()" onfocus="document.getElementById('work-attribution').select();" />
		  <input id="license-code" type="hidden" value="CC BY 3.0" />
		  <input id="license-url" type="hidden"
           value="http://creativecommons.org/licenses/by/3.0/hk/" />
		<a href="" id="attribution_help" class="helpLink">
		  <img src="http://creativecommons.org/@@/cc/images/information.png"
         alt="Information" />
		</a>
		</p>
		<div id="help_attribution_help" class="help_panel">
		  <div class="hd">
		    What does "Attribute this work" mean?
		  </div>
		  <div class="bd">
		    The page you came from contained embedded licensing
		    metadata, including how the creator wishes to be 
		    attributed for re-use.  You can use the HTML here to
		    cite the work.  Doing so will also include metadata on
		    your page so that others can find the original work as
		    well.
  		  </div>
		</div>

	      

            </li>

	  </ul>
	</div>
	<div id="deed-understanding">
	  <h3>With the understanding that:</h3>

	  <ul class="understanding license-properties">
            <li class="license">
	      <strong>Waiver</strong>
	      &mdash;
	      
		Any of the above conditions can be <a href="#" id="waived" class="helpLink">waived</a> if you get
		permission from the copyright holder.
	      
	    </li>
	      
	    <li class="license">
	      <strong>Other Rights</strong>
	      &mdash; 
	      In no way are any of the following rights affected by the license:
	     
	      <ul>

		<li>Your fair dealing
		  or <a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#Do_Creative_Commons_licenses_affect_fair_use.2C_fair_dealing_or_other_exceptions_to_copyright.3F" id="fair_use" class="helpLink">fair use</a> rights;
		</li>

		
		  <li>
		    The author's <a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#I_don.E2.80.99t_like_the_way_a_person_has_used_my_work_in_a_derivative_work_or_included_it_in_a_collective_work.3B_what_can_I_do.3F" id="moral_rights" class="helpLink">moral</a> rights;
		  </li>
		
		

		<li>
		  Rights other persons may have either in the work
		  itself or in how the work is used, such as 
		  <a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#When_are_publicity_rights_relevant.3F" id="publicity_rights" class="helpLink">publicity</a> or privacy rights.
		</li>
	      </ul>
	    </li>

            <li rel="cc:requires" resource="http://creativecommons.org/ns#Notice">
	      <strong>Notice</strong>
	      &mdash;
	      Vid all återanvändning och distribution måste du informera om licensvillkoren som gäller för verket. Det bästa sättet att göra detta är genom en länk till den här webbsidan.
	    </li>

          </ul>

          

          <div id="help_waived" class="help_panel">
            <div class="hd">What does "conditions can be waived" mean?</div>
            <div class="bd">
              <p>CC licenses anticipate that a licensor may want to
		waive compliance with a specific condition, such as
		attribution.</p>
              <p><a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#Can_I_change_the_terms_of_a_CC_license_or_waive_some_of_its_conditions.3F">Learn more</a>.</p>
            </div>
          </div>

          <div id="help_fair_use" class="help_panel">
            <div class="hd">What does "Fair use" mean?</div>
            <div class="bd">
              <p>All jurisdictions
              allow some limited uses of copyrighted material without
              permission.  CC licenses do not affect the rights of
              users under those copyright limitations and exceptions,
              such as fair use and fair dealing where applicable.</p>

              <p><a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#Do_Creative_Commons_licenses_affect_fair_use.2C_fair_dealing_or_other_exceptions_to_copyright.3F">Learn more</a>.</p>
            </div>
          </div>

          <div id="help_moral_rights" class="help_panel">
            <div class="hd">What are "Moral Rights"?</div>
            <div class="bd">
              <p>In addition to the right of licensors to request removal of their name from the work when used in a derivative or collective they don't like, copyright laws in most jurisdictions around the world (with the notable exception of the US except in very limited circumstances) grant creators "moral rights" which may provide some redress if a derivative work represents a "derogatory treatment" of the licensor's work.</p>

              <p><a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#I_don.E2.80.99t_like_the_way_a_person_has_used_my_work_in_a_derivative_work_or_included_it_in_a_collective_work.3B_what_can_I_do.3F">Learn more</a>.</p>

            </div>
          </div>

          <div id="help_publicity_rights" class="help_panel">
            <div class="hd">What are "Publicity Rights"?</div>
            <div class="bd">
              <p>Publicity
              rights allow individuals to control how their voice,
              image or likeness is used for commercial purposes in
              public.  If a CC-licensed work includes the voice or
              image of anyone other than the licensor, a user of the
              work may need to get permission from those individuals
              before using the work for commercial purposes.</p>

              <p><a href="http://wiki.creativecommons.org/Frequently_Asked_Questions#When_are_publicity_rights_relevant.3F">Learn more</a>.</p>
            </div>
          </div>
	  
        </div>
    <span id="referrer-metadata-container" />

       </div>
      </div>

      <div id="deed-foot">
        

          

	  
	    <a href="#" id="disclaimer" class="helpLink">Friskrivning</a>
	    <div id="help_disclaimer">
	      <div class="hd">Friskrivning</div>
	      <div class="bd"><p>
Commons Deed är inte en licens. Det är endast en enkel sammanfattning för att förstå licenstexten. Det är en lättläst version av några av de viktigaste villkoren. Se det som ett användarvänligt gränssnitt till Legal Code. Commons Deed har ingen juridisk relevans och dess innehåll återfinns inte i licenstexten.
</p>

<p>
Creative Commons är inte en advokatbyrå eller juridisk byrå och tillhandahåller inte juridiska tjänster. Att distribuera, visa eller länka till detta Commons Deed skapar inte ett klientförhållande.
</p></div>
	    </div>
	  

	<p style="text-align:center">

    

    

    

    Detta är en lättläst sammanfattning av <a href="legalcode" class="fulltext">licenstexten</a>.
 </p>

         
       </div>
    </div>
    <p id="footer">
      
      <a id="get_this"
         href="/license/results-one?license_code=by&amp;jurisdiction=hk&amp;version=3.0&amp;lang=sv">Use this license for your own work.</a>
      
    </p>

  </body>
</html>
