<html xmlns="http://www.w3.org/1999/xhtml"
      xmlns:cc="http://creativecommons.org/ns#"
      xmlns:dc="http://purl.org/dc/elements/1.1/">
  <head>
    <title>Creative Commons 
    Attribution-Noncommercial-No Derivative Works 2.5 Netherlands
  </title>

    <base href="http://creativecommons.org/licenses/by-nc-nd/2.5/nl/" /><link
    rel="stylesheet" type="text/css"
    href="http://creativecommons.org/licenses/@@/cc/includes/deed3.css"
    media="screen" />
    
    <link rel="stylesheet" type="text/css"
          href="http://creativecommons.org/licenses/@@/cc/includes/deed3-print.css"
          media="print" />

    <!--[if lt IE 7]><link rel="stylesheet" type="text/css" href="/includes/deed3-ie.css" media="screen" tal:attributes="href context/++resource++cc/includes/deed3-ie.css" /><![endif]-->

    <link rel="alternate" type="application/rdf+xml" href="rdf" /> 
    

<script type="text/javascript">
function setCookie(name, value, expires, path, domain, secure) {
    document.cookie= name + "=" + escape(value) +
        ((expires) ? "; expires=" + expires.toGMTString() : "") +
        ((path) ? "; path=" + path : "") +
        ((domain) ? "; domain=" + domain : "") +
        ((secure) ? "; secure" : "");
}
var expiry = new Date();
expiry.setTime(expiry.getTime()+(5*365*24*60*60*1000));
setCookie('lang','%s', expiry, '/');
</script>


    <script type="text/javascript"
            src="http://creativecommons.org/licenses/@@/cc/includes/referrer/ccdeed.js">
    </script>
    <script src="http://www.google-analytics.com/urchin.js" type="text/javascript"></script>
    <script type="text/javascript">
        _uacct="UA-2010376-1";  urchinTracker();
    </script>

   

  </head>
  <body onload="referrerMetadata()">

    <!-- 
<rdf:RDF xmlns="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <License rdf:about="http://creativecommons.org/licenses/by-nc-nd/2.5/nl/">
        <permits rdf:resource="http://creativecommons.org/ns#Reproduction"/>
        <permits rdf:resource="http://creativecommons.org/ns#Distribution"/>
        <requires rdf:resource="http://creativecommons.org/ns#Notice"/>
        <requires rdf:resource="http://creativecommons.org/ns#Attribution"/>
        <prohibits rdf:resource="http://creativecommons.org/ns#CommercialUse"/>
      </License>
    </rdf:RDF>
   -->

    <div id="header">
    <p align="center"><a href="/">Creative Commons</a></p>

    

<div style="width: 620px; margin-left: auto; margin-right: auto; text-align: center;">
<span align="left" dir="">This page is available in the following languages:</span>
<br />



<a href="./deed.af" title="Afrikaans" hreflang="af"
   rel="alternate nofollow" lang="af">Afrikaans</a>




<a href="./deed.bg" title="български" hreflang="bg"
   rel="alternate nofollow" lang="bg">български</a>




<a href="./deed.ca" title="Català" hreflang="ca"
   rel="alternate nofollow" lang="ca">Català</a>




<a href="./deed.da" title="Dansk" hreflang="da"
   rel="alternate nofollow" lang="da">Dansk</a>




<a href="./deed.de" title="Deutsch" hreflang="de"
   rel="alternate nofollow" lang="de">Deutsch</a>




<a href="./deed.en" title="English" hreflang="en"
   rel="alternate nofollow" lang="en">English</a>




<a href="./deed.en_CA" title="English (CA)" hreflang="en_CA"
   rel="alternate nofollow" lang="en_CA">English (CA)</a>




<a href="./deed.en_GB" title="English (GB)" hreflang="en_GB"
   rel="alternate nofollow" lang="en_GB">English (GB)</a>




<a href="./deed.en_US" title="English (US)" hreflang="en_US"
   rel="alternate nofollow" lang="en_US">English (US)</a>




<a href="./deed.eo" title="Esperanto" hreflang="eo"
   rel="alternate nofollow" lang="eo">Esperanto</a>




<a href="./deed.es" title="Castellano" hreflang="es"
   rel="alternate nofollow" lang="es">Castellano</a>




<a href="./deed.es_AR" title="Castellano (AR)"
   hreflang="es_AR" rel="alternate nofollow" lang="es_AR">Castellano (AR)</a>




<a href="./deed.es_CL" title="Español (CL)" hreflang="es_CL"
   rel="alternate nofollow" lang="es_CL">Español (CL)</a>




<a href="./deed.es_CO" title="Spanish (CO)" hreflang="es_CO"
   rel="alternate nofollow" lang="es_CO">Spanish (CO)</a>




<a href="./deed.es_MX" title="Castellano (MX)"
   hreflang="es_MX" rel="alternate nofollow" lang="es_MX">Castellano (MX)</a>




<a href="./deed.es_PE" title="Castellano (PE)"
   hreflang="es_PE" rel="alternate nofollow" lang="es_PE">Castellano (PE)</a>




<a href="./deed.eu" title="Euskara" hreflang="eu"
   rel="alternate nofollow" lang="eu">Euskara</a>




<a href="./deed.fi" title="Suomeksi" hreflang="fi"
   rel="alternate nofollow" lang="fi">Suomeksi</a>




<a href="./deed.fr" title="français" hreflang="fr"
   rel="alternate nofollow" lang="fr">français</a>




<a href="./deed.fr_CA" title="français (CA)"
   hreflang="fr_CA" rel="alternate nofollow" lang="fr_CA">français (CA)</a>




<a href="./deed.gl" title="Galego" hreflang="gl"
   rel="alternate nofollow" lang="gl">Galego</a>




<a href="./deed.he" title="עברית" hreflang="he"
   rel="alternate nofollow" lang="he">עברית</a>




<a href="./deed.hr" title="hrvatski" hreflang="hr"
   rel="alternate nofollow" lang="hr">hrvatski</a>




<a href="./deed.hu" title="Magyar" hreflang="hu"
   rel="alternate nofollow" lang="hu">Magyar</a>




<a href="./deed.it" title="Italiano" hreflang="it"
   rel="alternate nofollow" lang="it">Italiano</a>




<a href="./deed.ja" title="日本語" hreflang="ja"
   rel="alternate nofollow" lang="ja">日本語</a>




<a href="./deed.ko" title="한국어" hreflang="ko"
   rel="alternate nofollow" lang="ko">한국어</a>




<a href="./deed.mk" title="Macedonian" hreflang="mk"
   rel="alternate nofollow" lang="mk">Macedonian</a>




<a href="./deed.ms" title="Melayu" hreflang="ms"
   rel="alternate nofollow" lang="ms">Melayu</a>




<a href="./deed.nl" title="Nederlands" hreflang="nl"
   rel="alternate nofollow" lang="nl">Nederlands</a>




<a href="./deed.nso" title="Sesotho sa Leboa" hreflang="nso"
   rel="alternate nofollow" lang="nso">Sesotho sa Leboa</a>




<a href="./deed.pl" title="polski" hreflang="pl"
   rel="alternate nofollow" lang="pl">polski</a>




<a href="./deed.pt" title="Português" hreflang="pt"
   rel="alternate nofollow" lang="pt">Português</a>




<a href="./deed.sl" title="slovenski jezik" hreflang="sl"
   rel="alternate nofollow" lang="sl">slovenski jezik</a>




<a href="./deed.st" title="Sotho" hreflang="st"
   rel="alternate nofollow" lang="st">Sotho</a>




<a href="./deed.sv" title="svenska" hreflang="sv"
   rel="alternate nofollow" lang="sv">svenska</a>




<a href="./deed.zh" title="简体中文" hreflang="zh"
   rel="alternate nofollow" lang="zh">简体中文</a>




<a href="./deed.zh_TW" title="華語 (台灣)" hreflang="zh_TW"
   rel="alternate nofollow" lang="zh_TW">華語 (台灣)</a>




<a href="./deed.zu" title="isiZulu" hreflang="zu"
   rel="alternate nofollow" lang="zu">isiZulu</a>


</div>


    </div>

    <div id="deed" align="left" class="yellow" dir="">  
      <div id="deed-head">
	      <div id="cc-logo"><img src="/images/deed/cc-logo.jpg" alt="cc logo" /></div>
	      <h1><span>Creative Commons License Deed</span></h1>
        <div id="deed-license">
	        <h2 property="dc:title">Erkännande-Ickekommersiell-Inga bearbetningar 2.5 Nederländerna</h2>
        </div>
      </div>

      <div id="deed-main" align="left" dir="">
       <div id="deed-main-content">
          
        

        <div id="deed-rights" align="left" dir="">

        

<a href="/worldwide/nl/"><img
    src="/images/international/nl.png" border="0" /></a>
<h3 rel="cc:permits"
    href="http://creativecommons.org/ns#Reproduction">Du får:</h3>
		      <ul>
			<li class="license share" rel="cc:permits"
       href="http://creativecommons.org/ns#Distribution"><strong>att Dela</strong> — att kopiera, distribuera och sända verket</li>
			      
<span id="devnations-container" />
		      </ul>
        </div>
        <div id="deed-conditions">
		      <h3>På följande villkor:</h3>
	        <ul align="left" dir=""> 
            <li rel="cc:requires"
                href="http://creativecommons.org/ns#Attribution"
                class="license by">
	            <p><strong>Erkännande</strong>. 
              <span id="attribution-container">Du måste ange upphovsmannen och/eller licensgivaren på det sätt de anger (men inte på ett sätt som antyder att de godkänt eller rekommenderar din använding av verket).</span>
              
              <span id="by-more-container" /></p>
            </li>
            <li rel="cc:prohibits"
                href="http://creativecommons.org/ns#CommercialUse"
                class="license nc-eu">
	            <p><strong>Ickekommersiell</strong>. 
              
              <span>Du får inte använda verket för kommersiella ändamål.</span>
              <span id="nc-eu-more-container" /></p>
            </li>
            <li rel="" href="" class="license nd">
	            <p><strong>Inga bearbetningar</strong>. 
              
              <span>Du får inte förändra, bearbeta eller bygga vidare på verket.</span>
              <span id="nd-more-container" /></p>
            </li>
            <li id="more-container" class="license-hidden" />
            <li rel="cc:requires"
                href="http://creativecommons.org/ns#Notice">Vid all återanvändning och distribution måste du informera om licensvillkoren som gäller för verket. Det bästa sättet att göra detta är genom en länk till den här webbsidan.</li>
            <li>Undantag från villkoren ovan kan meddelas av upphovsrättsinnehavaren.</li>
            
            <li>Ingenting i denna licens begränsar upphovsmannens ideella rätt.</li>
            
            
          </ul>

          <div id="deed-newer">
    	      <p>Det finns en <a href="http://creativecommons.org/licenses/by-nc-nd/3.0/nl/">ny version</a> av denna licens. Du bör använda den för nya verk och överväga att omlicensiera existerande verk med den. Inga verk blir dock <em>automatiskt</em> licensierade under den nya licensen.</p>
          </div>

          </div>
    <span id="referrer-metadata-container" />

       </div>
      </div>


       <div id="deed-foot">
          

        
	<p id="disclaimer">
          <a href="/licenses/disclaimer-popup"
             onclick="window.open('/licenses/disclaimer-popup', 'characteristic_help', 'width=375,height=300,scrollbars=yes,resizable=yes,toolbar=no,directories=no,location=yes,menubar=no,status=yes'); return false;">Friskrivning</a> 
          <a href="/licenses/disclaimer-popup"
             onclick="window.open('/licenses/disclaimer-popup', 'characteristic_help', 'width=375,height=300,scrollbars=yes,resizable=yes,toolbar=no,directories=no,location=yes,menubar=no,status=yes'); return false;">
            <img src="/images/popup.gif" width="15" height="13" alt="disclaimer" border="0" /></a>
  	</p>
        <p align="center" style="margin-top:40px">
	  <strong>Dina lagstadgade rättigheter påverkas inte av denna licens.</strong>
	</p>

	<p align="center">

    

    

    

    Detta är en lättläst sammanfattning av <a href="legalcode" class="fulltext">licenstexten</a>.
 </p>

         
       </div>
    </div>
    <p id="footer">
      <a href="/about/licenses">Läs om hur du kan använda denna licens för dina verk</a>
    </p>

  </body>
</html>
