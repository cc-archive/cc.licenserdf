<html xmlns="http://www.w3.org/1999/xhtml"
      xmlns:cc="http://creativecommons.org/ns#"
      xmlns:dc="http://purl.org/dc/elements/1.1/">
  <head>
    <title>Creative Commons 
    Attribution 2.5 Canada
  </title>

    <!--<base href="" tal:attributes="href context/license/uri" />--><link rel="stylesheet" type="text/css" href="http://yui.yahooapis.com/2.5.1/build/container/assets/skins/sam/container.css" /> 

    <link rel="stylesheet" type="text/css"
          href="http://creativecommons.org/licenses/@@/cc/includes/deed3.css"
          media="screen" />
    
    <link rel="stylesheet" type="text/css"
          href="http://creativecommons.org/licenses/@@/cc/includes/deed3-print.css"
          media="print" />

    <!--[if lt IE 7]><link rel="stylesheet" type="text/css" href="/includes/deed3-ie.css" media="screen" tal:attributes="href context/++resource++cc/includes/deed3-ie.css" /><![endif]-->

    <link rel="alternate" type="application/rdf+xml" href="rdf" /> 
    

<script type="text/javascript">
function setCookie(name, value, expires, path, domain, secure) {
    document.cookie= name + "=" + escape(value) +
        ((expires) ? "; expires=" + expires.toGMTString() : "") +
        ((path) ? "; path=" + path : "") +
        ((domain) ? "; domain=" + domain : "") +
        ((secure) ? "; secure" : "");
}
var expiry = new Date();
expiry.setTime(expiry.getTime()+(5*365*24*60*60*1000));
setCookie('lang','%s', expiry, '/');
</script>



    <script type="text/javascript" src="http://yui.yahooapis.com/2.5.1/build/yahoo-dom-event/yahoo-dom-event.js">
    </script> 
    <script type="text/javascript" src="http://yui.yahooapis.com/2.5.1/build/connection/connection-min.js">
    </script> 
    <script type="text/javascript" src="http://yui.yahooapis.com/2.5.1/build/json/json-min.js">
    </script>

    <script type="text/javascript"
            src="http://creativecommons.org/licenses/@@/cc/includes/referrer/deed.js">
    </script>
    

    <script type="text/javascript" src="http://yui.yahooapis.com/2.5.1/build/container/container-min.js">
    </script>

    <script type="text/javascript"
            src="http://creativecommons.org/licenses/@@/cc/includes/deed3.js">
    </script>

    <script src="http://www.google-analytics.com/urchin.js" type="text/javascript"></script>
    <script type="text/javascript">
        _uacct="UA-2010376-1";  urchinTracker();
    </script>

   

  </head>
  <body class="yui-skin-sam">

    <!-- 
<rdf:RDF xmlns="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <License rdf:about="http://creativecommons.org/licenses/by/2.5/ca/">
        <permits rdf:resource="http://creativecommons.org/ns#Reproduction"/>
        <permits rdf:resource="http://creativecommons.org/ns#Distribution"/>
        <requires rdf:resource="http://creativecommons.org/ns#Notice"/>
        <requires rdf:resource="http://creativecommons.org/ns#Attribution"/>
        <permits rdf:resource="http://creativecommons.org/ns#DerivativeWorks"/>
      </License>
    </rdf:RDF>
   -->

    <div id="header">
    <p align="center">
      <a rel="dc:creator" href="http://creativecommons.org/">
	<span property="dc:title">Creative Commons</span>
    </a></p>

    

<div style="width: 620px; margin-left: auto; margin-right: auto; text-align: center;">
<span align="left" dir="">Denna sida finns tillgänglig på följande språk:</span>
<br />



<a href="./deed.af" title="Afrikaans" hreflang="af"
   rel="alternate nofollow" lang="af">Afrikaans</a>




<a href="./deed.bg" title="български" hreflang="bg"
   rel="alternate nofollow" lang="bg">български</a>




<a href="./deed.ca" title="Català" hreflang="ca"
   rel="alternate nofollow" lang="ca">Català</a>




<a href="./deed.da" title="Dansk" hreflang="da"
   rel="alternate nofollow" lang="da">Dansk</a>




<a href="./deed.de" title="Deutsch" hreflang="de"
   rel="alternate nofollow" lang="de">Deutsch</a>




<a href="./deed.el" title="Ελληνικά" hreflang="el"
   rel="alternate nofollow" lang="el">Ελληνικά</a>




<a href="./deed.en" title="English" hreflang="en"
   rel="alternate nofollow" lang="en">English</a>




<a href="./deed.en_CA" title="English (CA)" hreflang="en_CA"
   rel="alternate nofollow" lang="en_CA">English (CA)</a>




<a href="./deed.en_GB" title="English (GB)" hreflang="en_GB"
   rel="alternate nofollow" lang="en_GB">English (GB)</a>




<a href="./deed.en_US" title="English (US)" hreflang="en_US"
   rel="alternate nofollow" lang="en_US">English (US)</a>




<a href="./deed.eo" title="Esperanto" hreflang="eo"
   rel="alternate nofollow" lang="eo">Esperanto</a>




<a href="./deed.es" title="Castellano" hreflang="es"
   rel="alternate nofollow" lang="es">Castellano</a>




<a href="./deed.es_AR" title="Castellano (AR)"
   hreflang="es_AR" rel="alternate nofollow" lang="es_AR">Castellano (AR)</a>




<a href="./deed.es_CL" title="Español (CL)" hreflang="es_CL"
   rel="alternate nofollow" lang="es_CL">Español (CL)</a>




<a href="./deed.es_CO" title="Castellano (CO)"
   hreflang="es_CO" rel="alternate nofollow" lang="es_CO">Castellano (CO)</a>




<a href="./deed.es_EC" title="Español (Ecuador)"
   hreflang="es_EC" rel="alternate nofollow" lang="es_EC">Español (Ecuador)</a>




<a href="./deed.es_MX" title="Castellano (MX)"
   hreflang="es_MX" rel="alternate nofollow" lang="es_MX">Castellano (MX)</a>




<a href="./deed.es_PE" title="Castellano (PE)"
   hreflang="es_PE" rel="alternate nofollow" lang="es_PE">Castellano (PE)</a>




<a href="./deed.eu" title="Euskara" hreflang="eu"
   rel="alternate nofollow" lang="eu">Euskara</a>




<a href="./deed.fi" title="Suomeksi" hreflang="fi"
   rel="alternate nofollow" lang="fi">Suomeksi</a>




<a href="./deed.fr" title="français" hreflang="fr"
   rel="alternate nofollow" lang="fr">français</a>




<a href="./deed.fr_CA" title="français (CA)"
   hreflang="fr_CA" rel="alternate nofollow" lang="fr_CA">français (CA)</a>




<a href="./deed.gl" title="Galego" hreflang="gl"
   rel="alternate nofollow" lang="gl">Galego</a>




<a href="./deed.he" title="עברית" hreflang="he"
   rel="alternate nofollow" lang="he">עברית</a>




<a href="./deed.hr" title="hrvatski" hreflang="hr"
   rel="alternate nofollow" lang="hr">hrvatski</a>




<a href="./deed.hu" title="Magyar" hreflang="hu"
   rel="alternate nofollow" lang="hu">Magyar</a>




<a href="./deed.it" title="Italiano" hreflang="it"
   rel="alternate nofollow" lang="it">Italiano</a>




<a href="./deed.ja" title="日本語" hreflang="ja"
   rel="alternate nofollow" lang="ja">日本語</a>




<a href="./deed.ko" title="한국어" hreflang="ko"
   rel="alternate nofollow" lang="ko">한국어</a>




<a href="./deed.mk" title="Macedonian" hreflang="mk"
   rel="alternate nofollow" lang="mk">Macedonian</a>




<a href="./deed.ms" title="Melayu" hreflang="ms"
   rel="alternate nofollow" lang="ms">Melayu</a>




<a href="./deed.nl" title="Nederlands" hreflang="nl"
   rel="alternate nofollow" lang="nl">Nederlands</a>




<a href="./deed.nso" title="Sesotho sa Leboa" hreflang="nso"
   rel="alternate nofollow" lang="nso">Sesotho sa Leboa</a>




<a href="./deed.pl" title="polski" hreflang="pl"
   rel="alternate nofollow" lang="pl">polski</a>




<a href="./deed.pt" title="Português" hreflang="pt"
   rel="alternate nofollow" lang="pt">Português</a>




<a href="./deed.ro" title="română" hreflang="ro"
   rel="alternate nofollow" lang="ro">română</a>




<a href="./deed.sl" title="slovenski jezik" hreflang="sl"
   rel="alternate nofollow" lang="sl">slovenski jezik</a>




<a href="./deed.sr" title="српски " hreflang="sr"
   rel="alternate nofollow" lang="sr">српски </a>




<a href="./deed.sr_LATN" title="srpski (latinica)"
   hreflang="sr_LATN" rel="alternate nofollow"
   lang="sr_LATN">srpski (latinica)</a>




<a href="./deed.st" title="Sotho" hreflang="st"
   rel="alternate nofollow" lang="st">Sotho</a>




<a href="./deed.sv" title="svenska" hreflang="sv"
   rel="alternate nofollow" lang="sv">svenska</a>




<a href="./deed.zh" title="中文" hreflang="zh"
   rel="alternate nofollow" lang="zh">中文</a>




<a href="./deed.zh_TW" title="華語 (台灣)" hreflang="zh_TW"
   rel="alternate nofollow" lang="zh_TW">華語 (台灣)</a>




<a href="./deed.zu" title="isiZulu" hreflang="zu"
   rel="alternate nofollow" lang="zu">isiZulu</a>


</div>


    </div>

    <div id="deed" align="left" class="green" dir="">  
      <div id="deed-head">
	      <div id="cc-logo"><img src="/images/deed/cc-logo.jpg" alt="cc logo" /></div>
	      <h1><span>Creative Commons License Deed</span></h1>
        <div id="deed-license">
	        <h2 property="dc:title">Erkännande 2.5 Kanada</h2>
        </div>
      </div>

      <div id="deed-main" align="left" dir="">
       <div id="deed-main-content">
          
  <div id="libre">
    <a href="http://freedomdefined.org/">
      <img src="/images/deed/seal.png" border="0"
           alt="This license is acceptable for Free Cultural Works." />
    </a>
  </div>

        <div id="deed-rights" align="left" dir="">

        

<a href="/worldwide/ca/"><img
    src="/images/international/ca.png" border="0" /></a>
<h3 rel="cc:permits"
    href="http://creativecommons.org/ns#Reproduction">Du får:</h3>
		      <ul>
			<li class="license share" rel="cc:permits"
       href="http://creativecommons.org/ns#Distribution"><strong>att Dela</strong> — att kopiera, distribuera och sända verket</li>
			      <li class="license remix" rel="cc:permits"
             href="http://creativecommons.org/ns#DerivativeWorks"><strong>att Remixa</strong> — att skapa bearbetningar</li>
            <li id="more-container" class="license-hidden" />
	    <span id="devnations-container" />
		      </ul>
        </div>
        <div id="deed-conditions">
	  <h3>På följande villkor:</h3>

	  <ul align="left" dir=""> 
            <li rel="cc:requires"
                href="http://creativecommons.org/ns#Attribution"
                class="license by">
	      <p><strong>Erkännande</strong>. 
		<span id="attribution-container">Du måste ange upphovsmannen och/eller licensgivaren på det sätt de anger (men inte på ett sätt som antyder att de godkänt eller rekommenderar din använding av verket).</span>
		
		<span id="by-more-container" />
	      </p>

	      
		<p id="work-attribution-container" style="display:none;">
		  <strong>Attribute this work:</strong><br />
		  <input id="work-attribution" value="" type="text" readonly onclick="this.select()" onfocus="document.getElementById('work-attribution').select();" />
		  <input id="license-code" type="hidden" value="CC BY 2.5" />
		  <input id="license-url" type="hidden"
           value="http://creativecommons.org/licenses/by/2.5/ca/" />
		<a href="" id="attribution_help">
		  <img src="http://creativecommons.org/licenses/@@/cc/images/information.png" />
		</a>
		</p>
		<div id="attribution_help_panel">
		  <div class="hd">
		    What does "Attribute this work" mean?
		  </div>
		  <div class="bd">
		    The page you came from contained embedded licensing
		    metadata, including how the creator wishes to be 
		    attributed for re-use.  You can use the HTML here to
		    cite the work.  Doing so will also include metadata on
		    your page so that others can find the original work as
		    well.
  		  </div>
		</div>

	      

            </li>
            <li rel="cc:requires"
                href="http://creativecommons.org/ns#Notice">Vid all återanvändning och distribution måste du informera om licensvillkoren som gäller för verket. Det bästa sättet att göra detta är genom en länk till den här webbsidan.</li>
            <li>Undantag från villkoren ovan kan meddelas av upphovsrättsinnehavaren.</li>
            
            <li>Ingenting i denna licens begränsar upphovsmannens ideella rätt.</li>
            
            
          </ul>

          

          </div>
    <span id="referrer-metadata-container" />

       </div>
      </div>


      <div id="deed-foot">
        

          

	  
	    <a href="" id="disclaimer">Friskrivning</a>
	    <div id="disclaimer_panel">
	      <div class="hd">Friskrivning</div>
	      <div class="bd"><p>
Commons Deed är inte en licens. Det är endast en enkel sammanfattning för att förstå licenstexten. Det är en lättläst version av några av de viktigaste villkoren. Se det som ett användarvänligt gränssnitt till Legal Code. Commons Deed har ingen juridisk relevans och dess innehåll återfinns inte i licenstexten.
</p>

<p>
Creative Commons är inte en advokatbyrå eller juridisk byrå och tillhandahåller inte juridiska tjänster. Att distribuera, visa eller länka till detta Commons Deed skapar inte ett klientförhållande.
</p></div>
	  </div>
	  

        <p align="center" style="margin-top:40px">
	  <strong>Dina lagstadgade rättigheter påverkas inte av denna licens.</strong>
	</p>

	<p align="center">

    
     Detta är en lättläst sammanfattning av licenstexten som finns tillgänglig på följande språk:
       <br />

     

     
         <a href="legalcode.en">engelska</a> 
         <a href="legalcode.fr">franska</a>
     

     

     

     
    

    

    

    
 </p>

         
       </div>
    </div>
    <p id="footer">
      <a href="/about/licenses">Läs om hur du kan använda denna licens för dina verk</a>
    </p>

  </body>
</html>
